module led (
  input wire key_in,
  output wire key_out
);

assign key_out=key_in;

endmodule